`ifndef BOARD_PKG_SVH
`define BOARD_PKG_SVH

package board_pkg;

    parameter KEYS_W    = 3;
    parameter LEDS_W    = 2;
    parameter VGA_RGB_W = 3;

endpackage : board_pkg

`endif 
