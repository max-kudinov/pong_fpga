(* blackbox *)
module TLVDS_OBUF (I, O, OB);
  input I;
  output O;
  output OB;
endmodule

