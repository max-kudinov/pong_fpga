`ifndef LFSR_PKG_SVHH
`define LFSR_PKG_SVHH

package lfsr_pkg;

    parameter RND_NUM_W = 9;
    parameter RND_SEED  = 1337;
    parameter TAPS      = 'h110;

endpackage : lfsr_pkg

`endif
