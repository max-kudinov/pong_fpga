`include "sprite_pkg.svh"

interface sprite_if;
    import sprite_pkg::sprite_t;

    sprite_t sprite;

endinterface : sprite_if
